Caleb Alexander
vi 1 0 ac 1

R1 2 1 22.85k
R2 3 2 1.273k

C1 3 0 1.5n
C2 4 2 15n

X1 3 4 4 OPAMP


*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP

.AC DEC 100 100 100K
.PROBE
.END