Caleb Alexander
vi 1 0 ac 1
R3 2 0 212
R2 3 2 212
R1 4 3 1.7k
C1 4 3 0.015uF
X1 1 2 4 OPAMP
*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP
.AC DEC 100 100 100K
.PROBE
.END
