Caleb Alexander
vi 1 0 ac 1

C1 2 1 15n
C2 3 2 15n

R1 3 0 1.7k
R2 4 2 1.7k

X1 3 4 4 OPAMP


*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP

.AC DEC 100 100 100K
.PROBE
.END