Caleb Alexander
vi 1 0 ac 1
R1 2 1 425
R2 3 2 1.7k
C1 3 2 0.015uF
R3 4 3 4.25k
X1 0 3 4 OPAMP
*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP
.AC DEC 100 100 100K
.PROBE
.END
