Caleb Alexander
vi 1 0 ac 1
R1 3 1 1.7k
C1 2 1 0.015uF
R2 2 0 1.7k
R3 4 3 1.7k
X1 2 3 4 OPAMP
*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP
.AC DEC 100 100 100K
.PROBE
.END
