Caleb Alexander
vi 1 0 ac 1

R6 2 0 5.118k
C2 2 1 15n

R4 3 2 1.7k

C1 4 3 15n

R1 5 4 1.7k

R2 6 5 1.7k

R7 6 1 1.7k

X1 2 4 5 OPAMP
X2 6 4 3 OPAMP

*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP

.AC DEC 100 100 100K
.PROBE
.END