Caleb Alexander
vi 1 0 ac 1

R5 2 1 10.2k
R6 2 0 10.2k
C3 2 0 15n

R4 3 2 1.7k

C1 4 3 15n

R1 5 4 1.7k

R2 6 5 1.7k

R3 6 0 1.7k

X1 2 4 5 OPAMP
X2 6 4 3 OPAMP

*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP

.AC DEC 100 100 100K
.PROBE
.END