Caleb Alexander
VS	1	0	AC	1

C1	2	1	0.1u
R1	3	2	16k
C2	4	3	47p
R2	4	3	115k

XOP	0 3	4	OPAMP1


* OPAMP MACRO MODEL

.SUBCKT OPAMP1 1 2 3
RIN 1 2 2E6
GM1 4 0 1 2 1.38E-4
R3 4 0 1E5
CC 4 5 20E-12
GM2 5 0 4 0 106
R01 3 5 150
R02 5 0 150
.ENDS OPAMP1

* ANALYSIS
* .TRAN	0.1US	10US
.ac dec 2000 10 300000
.PROBE
.END
