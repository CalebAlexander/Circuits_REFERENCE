Caleb Alexander
vi 1 0 ac 1
R1 1 2 12k
R2 2 3 15k
R3 3 0 4.3k
C  2 3 22n
.ac dec 10 10 100000k
.probe
.end