Caleb Alexander
vi 1 0 PWL(0 10 3M 10)
R1 1 2 12k
R2 2 3 15k
R3 3 0 4.3k
C1 2 3 0.022u IC = 0
.tran 0 3M UIC
.probe
.end
