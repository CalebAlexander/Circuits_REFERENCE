Caleb Alexander
vi 1 0 PULSE(0 10 1p)
R1 1 2 68k
R2 2 0 33k
R3 2 3 6.8k
L1 3 4 3m
C1 4 0 1p
.tran 1n 2u
.print tran I(L1)
.end
