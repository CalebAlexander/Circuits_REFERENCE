Caleb Alexander
VI 1 0 AC 1 SIN(0 0.7 1K)
*VOLTAGE SOURCE FOR EITHER AC OR TRAN ANALYSIS, ARGUMENTS OF SINE DC LEVEL, AMPLITUDE, FREQ
RB1 2 0 73K
RB2 6 2 173K
RE1 4 0 4.3K
RE2 4 7 73
RC 6 3 7.3K
RL 5 0 4.3K
C1 1 2 0.22U
C2 3 5 10U
CE 7 0 100U
Q 3 2 4 QKITTYCAT
VPLUS 6 0 DC 15
.MODEL QKITTYCAT NPN(IS=6.734F BF=416 VA=74.03 CJC=3.638P TF=0.3012N RB=10)
*IS SATURATION CURRENT, BF FORWARD BETA, VA EARLY VOLTAGE,
*CJC COLLECTION JUNCTION CAPACITANCE, TF FORWARD TRANSIT TIME,
*RB BASE SPREADING RESISTANCE
*DO ONE ANALYSIS AT A TIME. PUT AN ASTERISK IN FRONT OF THE OTHERS
.OP
*OP PROVIDES THE Q POINT
*.AC DEC 300 10 100MEG
*.TRAN 0 3M
*.FOUR 1K V(5)
*FOURIER ANALYSIS OF VOLTAGE AT NODE 5 WITH 1K AS FUNDAMENTAL FREQUENCY
.PROBE
.END
