Caleb Alexander
vi 1 0 ac 1
C1 2 1 0.1uF
R1 2 0 255
R3 3 0 3k
R4 4 3 27k
X1 2 3 4 OPAMP
*QUASI-IDEAL OP-AMP SUBCIRCUIT
.SUBCKT OPAMP 1 2 3
EOUT 3 0 1 2 200K
.ENDS OPAMP
.AC DEC 100 100 100K
.PROBE
.END
