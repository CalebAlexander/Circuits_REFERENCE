Quadrature Oscillator
*With Diode Amplitude Limiter
R1 1 Vout1 2.5k
R2 3 Vout2 4.9k
R3 0 5 1k
R4 5 Vout1 1k
R5 3 Vout1 4k

VCC vcc 0 15
VEE vee 0 -15

R6 vee 6 30k
R7 vcc 2 30k
R8 Vout2 2 5.1k
R9 Vout2 6 5.1k

C1 1 Vout2 10n
C2 3 0 10n

D1 6 1 d1n4148
D2 1 2 d1n4148

X1 0 1 vcc vee Vout2 TL071
X2 3 5 vcc vee Vout1 TL071

.model d1n4148 D(is=1n bv=100 n=1.8)
* TL071 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.01 ON 06/16/89 AT 13:08
* (REV N/A) SUPPLY VOLTAGE: +/-15V
* CONNECTIONS: NON-INVERTING INPUT
* | INVERTING INPUT
* | | POSITIVE POWER SUPPLY
* | | | NEGATIVE POWER SUPPLY
* | | | | OUTPUT
* | | | | |
.SUBCKT TL071 1 2 3 4 5
*
C1 11 12 3.498E-12
C2 6 7 15.00E-12
DC 5 53 DX
DE 54 5 DX
DLP 90 91 DX
DLN 92 90 DX
DP 4 3 DX
EGND 99 0 POLY(2) (3,0) (4,0) 0 .5 .5
FB 7 99 POLY(5) VB VC VE VLP VLN 0 4.715E6 -5E6 5E6 5E6 -5E6
GA 6 0 11 12 282.8E-6
GCM 0 6 10 99 8.942E-9
ISS 3 10 DC 195.0E-6
HLIM 90 0 VLIM 1K
J1 11 2 10 JX
J2 12 1 10 JX
R2 6 9 100.0E3
RD1 4 11 3.536E3
RD2 4 12 3.536E3
RO1 8 5 150
RO2 7 99 150
RP 3 4 2.143E3
RSS 10 99 1.026E6
VB 9 0 DC 0
VC 3 53 DC 2.200
VE 54 4 DC 2.200
VLIM 7 8 DC 0
VLP 91 0 DC 25
VLN 0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=15.00E-12 BETA=270.1E-6 VTO=-1)
.ENDS TL071
.TRAN 0 8m UIC
.PROBE
