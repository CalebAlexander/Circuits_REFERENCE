Caleb Alexander
VS	1	0	AC	1

C1	2	0	0.1u
R1	3	2	53
R2	4	3	332

XOP	1 3	4	OPAMP2


* OPAMP MACRO MODEL

.SUBCKT OPAMP2 1 2 3
EOUT 3 0 1 2 300K
.ENDS OPAMP2

* ANALYSIS
* .TRAN	0.1US	10US
.ac dec 2000 10 300000
.PROBE
.END
